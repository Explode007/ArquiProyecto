module ConditionHandler(
    input B_in,
    input BL_in,
    input I_Cond_in,
    input Flags_in,

    output reg TA_Ctrl_out,
    output reg BL_COND_out,
    output reg COND_EVAL_out
);

endmodule