`include "Adder.v"
`include "ControlUnit.v"
`include "cuMux.v"
`include "PC.v"
`include "rom.v"
`include "fase3pipereg.v"

module PPU();

reg rst;
reg clk;
reg s;
//Wires & More!

//Preload
integer fi, code, i;
reg [7:0] data;
reg [8:0] Address;

//PC Wires
wire [31:0] PC_Out; 
wire [31:0] PC_In; 
reg LE;
wire [31:0] Adder_Out;

//ROM Wires
wire [31:0] insMem_Out;

//IF-ID Reg Wires
wire [11:0] imm_in;
wire [31:0] cu_in;

//Control Unit Wires
wire rf_en;
wire [3:0] alu_op;
wire Load;
wire branch_link;
wire s_bit;
wire rw;
wire size;
wire datamem_en;

//Control Unit Mux Wires
wire rf_en_out;
wire [3:0] alu_op_out;
wire Load_out;
wire branch_link_out;
wire s_bit_out;
wire rw_out;
wire size_out;
wire datamem_en_out;

//Instantiations here!
PC PCReg(
    .E(LE), 
    .Reset(rst), 
    .clk(clk), 
    .PC_In(PC_In), 
    .PC_Out(PC_Out)
);

adder add(
    .Adder_OUT(Adder_Out),
    .Adder_IN(PC_Out)
);

rom insMem(
    .I(insMem_Out),
    .A(PC_Out[7:0])
);

control_unit CU(
    .instruction(cu_in),
    .rf_en(rf_en),
    .alu_op(alu_op),
    .Load(Load),
    .branch_link(branch_link),
    .s_bit(s_bit),
    .rw(rw),
    .size(size),
    .datamem_en(datamem_en)
);

cuMux Mux(
    .s(s),
    .rf_en_in(rf_en),
    .alu_op_in(alu_op),
    .Load_in(Load),
    .branch_link_in(branch_link),
    .s_bit_in(s_bit),
    .rw_in(rw),
    .size_in(size),
    .datamem_en_in(datamem_en),

    .rf_en_out(rf_en_out),
    .alu_op_out(alu_op_out),
    .Load_out(Load_out),
    .branch_link_out(branch_link_out),
    .s_bit_out(s_bit_out),
    .rw_out(rw_out),
    .size_out(size_out),
    .datamem_en_out(datamem_en_out)
);

if_id_reg IF_ID(
    .clk(clk),
    .load_enable(LE),
    .reset(rst),

    .instruction(PC_Out),
    
    .cu_in(cu_in)
);

id_exe_reg ID_EXE(
    .clk(clk), 
    .reset(rst),

    .am,
    .alu_op,
    .rf_en,
    .s,
    .datamem_en,
    .readwrite,
    .size,
    .load_instruction,

    .am_out,
    .alu_op_out,
    .rf_en_out,
    .s_out,
    .datamem_en_out,
    .readwrite_out,
    .size_out,
    .load_instruction_out
);

exe_mem_reg EXE_MEM(
    .clk(clk),
    .reset(rst),

    .rf_en,
    .datamem_en,
    .readwrite,
    .size,
    .load_instruction,
    
    .rf_en_out,
    .datamem_en_out,
    .readwrite_out,
    .size_out,
    .load_instruction_out
);

mem_wb_reg MEM_WB(
    .clk(clk),
    .reset(rst),

    .rf_en,
    
    .rf_en_out
);

//Simulation stuff here!

initial begin
    fi = $fopen("testcode_Fase_III(2).txt","r");
    Address = 9'b000000000;
    while (!$feof(fi)) begin
        code = $fscanf(fi, "%b", data);
        insMem.Mem[Address] = data;
        Address = Address + 1;
    end
    $fclose(fi);
    
    LE = 1'b1;
    clk = 0;
    forever #2 clk = ~clk;
    rst = 1'b1;
    #3 rst = 1'b0;

    s = 1'b0;
    #32 s = 1'b1;

    $monitor("Time: %0t", 
    $time
    );
end

endmodule